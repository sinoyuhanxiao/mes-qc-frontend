VITE_API_URL=http://10.10.60.209:8090
VITE_QC_SUMMARY_API=http://10.10.60.209:8010
